-- Elementos de Sistemas
-- by Luciano Soares
-- FullAdder.vhd

-- Implementa Full Adder

Library ieee;
use ieee.std_logic_1164.all;

entity FullAdder is
	port(
		a,b,c:      in STD_LOGIC;   -- entradas
		soma,vaium: out STD_LOGIC   -- sum e carry
	);
end entity;

architecture rtl of FullAdder is

begin
<<<<<<< HEAD
	soma <= a xor b xor c;
	vaium <= (a and b) or (c and a) or (c and b);
=======

>>>>>>> upstream/master
end architecture;
